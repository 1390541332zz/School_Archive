/*---------------------------------------------------------------------------*
 * Module: Gameboy Memory Map Master                                         *
 * Purpose: Connects the Gameboy DMG to all memory mapped object: SD Card,   *
 *     Static DRAM, and DAC/VGA Configuration.                               *
 * Last Edit: 2019-04-30                                                     *
 * Maintainer: Jacob Abel                                                    *
 *---------------------------------------------------------------------------*/

module mm_cntrlr(
/*---------------------------------------------------------------------------*/
/*                                Variables                                  */
/*---------------------------------------------------------------------------*/
    mm_ebab.master mm
);

endmodule : mm_cntrlr
