module question4 (
    input [7:0] in,
    output [31:0] out );//


endmodule