module i2cmasterwrite(input      clk,
                      input  reset,
                      input  init,
                      output sck,
                      inout  sda
                      );
   

	// YOU HAVE TO DEVELOP THIS CODE
    // YOU ARE ALLOWED (AND ENCOURAGED) TO INTRODUCE NEW FILES, NEW MODULES
	// USE A HIERARCHICAL FSM, WITH BITXMIT THE FRONT-END
   
endmodule
