module question5 ( input clk, input reset, input d, output q );

endmodule

module my_dff ( input clk, input reset, input d, output reg q );


endmodule