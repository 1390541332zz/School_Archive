///Help
