// NAME YOUR MODULE TO REFLECT YOUR OWN PID.
// CHANGE THE INFORMATION IN THE HEADER BLOCK.
// SAVE THE FILE USING THE NEW FILE NAME. REMEMBER TO UPDATE YOUR PROJECT WITH THE RENAMED FILE.
// DELETE THESE COMMENTS AFTER YOU HAVE DONE THESE THINGS.

////////////////////////////////////////////////////////////////////////////////////////////////////
// Filename:    game_gate_YOURPID.v
// Author:   
// Date:        04 September 2018
// Version:     1
// Description: This is a structural model for the circuit that implements Project 1.
//              The circuit uses the inputs to determine which of two players, if either,
//              has won the game.

module game_gate_YOURPID(player_a, player_b, player_a_wins, player_b_wins, tie_game);
   input [1:0] player_a, player_b;
   output      player_a_wins, player_b_wins, tie_game;

   // YOU MAY DECLARE WIRES AS NEEDED.

   // INSERT YOUR CODE HERE.
    
endmodule
