module question6 ( 
    input clk,
	input reset,
    input [7:0] d, 
    input [1:0] sel, 
    output [7:0] q 
);

endmodule

module my_dff8 ( input clk, input reset, input [7:0] d, output reg [7:0] q );

endmodule