// synthesis verilog_input_version verilog_2001
module question10 (
    input [3:0] in,
    output reg [1:0] pos  );
    

endmodule