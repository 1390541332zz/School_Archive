////////////////////////////////////////////////////////////////////////////////////////////////////
// File: ECE2504SimpleComputer.v
// Top-level file for Simple Computer projects (Project 3, Project 4)
// The Simple Computer from Chapter 8
//
// ******************************************
// YOU ARE NOT PERMITTED TO MODIFY THIS FILE.
// ******************************************
//
// This is a simplified version of the simple computer module created by Xin Xin in June 2012.
//
// Created by Tom Martin, 11/29/2012
// Modified by P. Athanas, 3/2013
// Modified by KLC, 11/2013
// Modified by Hsiao, 10/2015
// Modified by KLC, 11/2015
//
// Changes:
// 1. The accelerometer has been removed.
// 2. The modules have been re-arranged in the files to indicate which modules can be changed and
//    which must not be changed.
// 3. This version uses all four DIP switches to control the LEDs instead of having one control
//    whether the clock is enabled by the pushbutton.
// 4. KEY0 is the reset and KEY1 is the clock enable to be consistent with Project 2.
// 5. The synthesis keep directive has been added to signals of interest in the cpu module.
// 6. Add toggling of LEDS using KEY[0] for SW[3:1] = 110 and 111 so that r6 and r7 can be
//    displayed. This might lead to poor behavior, but the board is input-constrained.
//
// ================================================
// This code is generated by Terasic System Builder
// ================================================
////////////////////////////////////////////////////////////////////////////////////////////////////

`timescale 1 ns/1 ps

module ECE2504SimpleComputer(CLOCK_50, KEY, SW, LED);

//=======================================================
//  PORT declarations
//=======================================================

	//////////// CLOCK //////////
	input        CLOCK_50;

	//////////// KEY //////////
	input [1:0]  KEY;

	//////////// SW //////////
	input [3:0]  SW;

	//////////// LED //////////
	output [7:0] LED;

//=======================================================
//  WIRE and REG declarations
//=======================================================

	wire        rst_inv;
	wire        cpu_clk;
	wire        cpu0_clk;
	wire        cpu0_clk_en;
	wire [15:0] r0, r1, r2, r3, r4, r5, r6, r7, IR, PC, mux6, mux7;
	reg         cpu0_clk_en_delay0, cpu0_clk_en_delay1;

//=======================================================
//  Structural coding
//=======================================================

	assign rst_inv = ~KEY[0]; // In this sense, rst_inv is an active low signal.
	assign cpu_clk = cpu0_clk;

	// Instantiate CPU.
	cpu cpu0
	(
		.rst(rst_inv),
		.clk(cpu_clk),
		.r0(r0),
		.r1(r1),
		.r2(r2),
		.r3(r3),
		.r4(r4),
		.r5(r5),
		.r6(r6),
		.r7(r7),
		.IR(IR),
		.PC(PC)
	);

	// Instantiate push-button finite state machine.
	// The FSM and clock assignments allow the CPU to use KEY1 as the clock signal. KEY1 is gated
	// with the 50 MHz clock to generate one 50 MHz clock pulse each time KEY1 is pushed. The FSM
	// generates one clock enable signal per button push.

	button_fsm button_fsm0
	(
		.rst(rst_inv),
		.clk(CLOCK_50),
		.button(KEY[1]),
		.cpu0_clk_en(cpu0_clk_en)
	);

	// This is Altera's recommended way to implement clock gating.

	always@(posedge CLOCK_50) //make sure cpu0_clk_en_delay0 is one clock cycle
		cpu0_clk_en_delay0 = cpu0_clk_en;

	always@(negedge CLOCK_50)
		cpu0_clk_en_delay1 = cpu0_clk_en_delay0;

	assign cpu0_clk = cpu0_clk_en_delay1 & CLOCK_50;

	// End of clock generation portion.

	// Use KEY[0] to select between PC/r6 and IR/r7 for LED display
	// When resetting the device (with KEY0 pressed), the PC will not be displayed, r6 will be.

	assign mux6 = KEY[0] ? PC : r6;
	assign mux7 = KEY[0] ? IR : r7;

	// Assign the LEDs based upon the DIP switch settings.

	mux16_1_8bits LED_mux(LED, SW, mux7[15:8], mux7[7:0], mux6[15:8], mux6[7:0], r5[15:8], r5[7:0], r4[15:8], r4[7:0],
                                  	r3[15:8],   r3[7:0],   r2[15:8],   r2[7:0], r1[15:8], r1[7:0], r0[15:8], r0[7:0]);

endmodule
