module question8(
    input [31:0] a,
    input [31:0] b,
    input sub,
    output [31:0] result
);

endmodule

module add1 ( input a, input b, input cin,   output sum, output cout );

endmodule

module add16 ( input[15:0] a, input[15:0] b, input cin, output[15:0] sum, output cout );

endmodule

